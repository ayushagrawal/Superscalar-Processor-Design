library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.components.all;

entity lst_unit is

		port(clk : in std_logic;
			  reset : in std_logic;
			  input : in std_logic_vector(42 downto 0);
			  output : out std_logic_vector(21 downto 0));
			  
end entity;

architecture lst_arch of lst_unit is
	
	
	
begin
	

	
end architecture;